module myand(y, a, b);
input a,b;
output y; 
  
//assign y=a&b;
and A1(y,a,b);
endmodule

