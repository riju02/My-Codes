module mynot(y, a);
input a;
output y; 
  
not A1(y,a);
endmodule

