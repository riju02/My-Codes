module myor(y, a,b);
input a,b;
output y; 
  
  or a2(y,a,b);
endmodule