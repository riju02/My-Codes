module mynot(y, a);
input a;
output y; 
  
//assign y=a&b;
not A1(y,a);
endmodule

